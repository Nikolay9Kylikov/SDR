`timescale 1ns/1ps

module cordic (
	input	clk_i,
	input	rst_i,
	input	valid_i,
	input	[31:0] phase_i,
	output	reg signed [15:0] sin_o,
	output	reg signed [15:0] cos_o,
	output	reg valid_o
);
	localparam [31:0] HALF_PI_PHASE = 32'h4000_0000; // 2^30 == π/2
	localparam [31:0] ATAN_TABLE [15:0] = {
		32'h0000517D, // i=15 (LS in this listing)  -- trimmed if ITER < 16
		32'h0000A2FA, // i=14
		32'h000145F3, // i=13
		32'h00028BE6, // i=12
		32'h000517CC, // i=11
		32'h000A2F98, // i=10
		32'h00145F2F, // i=9
		32'h0028BE53, // i=8
		32'h00517C55, // i=7
		32'h00A2F61E, // i=6
		32'h0145D7E1, // i=5
		32'h028B0D43, // i=4
		32'h051111D4, // i=3
		32'h09FB385B, // i=2
		32'h12E4051E, // i=1
		32'h20000000  // i=0  = pi/4 in phase units
	};

	reg signed [47:0] x_init;
	reg signed [47:0] y_init;
	reg signed [31:0] theta_init;
	
	reg [16:0] valid_stage;
	reg [33:0] quadrant;

	always @(posedge clk_i) begin
		if (rst_i) begin
			x_init <= 0;
			y_init <= 0;
			theta_init <= 32'sd0;
		end
		else begin
			valid_stage <= {valid_stage[15:0], valid_i};
			quadrant <= {quadrant[31:0], phase_i[31:30]};
			if (valid_i) begin
				x_init <= {16'b0, 32'h69648523}; // Q2.30 all numbers, because theta belongs [2pi:2pi]
				y_init <= 0;
				case(phase_i[31:30])
					2'b00: theta_init <= $signed({2'b0, phase_i[29:0]});								// 0..+pi/2
					2'b01: theta_init <= $signed(HALF_PI_PHASE) - $signed({2'b0, phase_i[29:0]});		// +pi/2 .. 0
					2'b10: theta_init <= $signed({2'b0, phase_i[29:0]});								// 0 .. -pi/2
					2'b11: theta_init <= -($signed(HALF_PI_PHASE) - $signed({2'b0, phase_i[29:0]}));	// -pi/2 .. 0
					default: theta_init <= 32'sd0;
				endcase
			end
			else begin
				x_init <= 0;
				y_init <= 0;
				theta_init <= 32'sd0;
			end
		end
	end

	reg signed [47:0] x [16:0]; //16 - number of iterations
	reg signed [47:0] y [16:0];
	reg signed [31:0] theta [16:0];

	always @(posedge clk_i) begin
		x[0]<= x_init;
		y[0]<= y_init;
		theta[0]<= theta_init;
	end

	genvar i;
	generate
		for (i = 0; i < 16; i = i + 1) begin : cordic_stages
			always @(posedge clk_i) begin
				if (rst_i) begin
					x[i+1] <= 0;
					y[i+1] <= 0;
					theta[i+1] <= 32'sd0;
				end
				else begin
					if (valid_stage[i]) begin
						if (theta[i] >= 0) begin
							x[i+1] <= x[i] - (y[i] >>> i);
							y[i+1] <= y[i] + (x[i] >>> i);
							theta[i+1] <= theta[i] - $signed(ATAN_TABLE[i]);
						end
						else begin
							x[i+1] <= x[i] + (y[i] >>> i);
							y[i+1] <= y[i] - (x[i] >>> i);
							theta[i+1] <= theta[i] + $signed(ATAN_TABLE[i]);
						end
					end
					else begin
						x[i+1]<= 0;
						y[i+1]<= 0;
						theta[i+1]<= 32'sd0;
					end
				end
			end
		end
	endgenerate
	
	always @(posedge clk_i) begin
		if (rst_i) begin
			valid_o <= 1'b0;
			cos_out <= 16'sd0;
			sin_out <= 16'sd0;
		end
		else begin
			valid_o <= valid_stage[16];
			case(quadrant[33:32])
				2'b00: begin
					cos_o <= $signed(x[16] >>> 32'd15);
					sin_o <= $signed(y[16] >>> 32'd15);
				end
				2'b01: begin
					cos_o <= -$signed(y[16] >>> 32'd15); 
					sin_o <= $signed(x[16] >>> 32'd15);
				end
				2'b10: begin
					cos_o <= -$signed(x[16] >>> 32'd15);
					sin_o <= -$signed(y[16] >>> 32'd15);
				end
				2'b11: begin
					cos_o <= -$signed(y[16] >>> 32'd15);
					sin_o <= -$signed(x[16] >>> 32'd15);
				end
			endcase
		end
	end

endmodule